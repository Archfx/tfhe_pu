`timescale 1 ps / 1 ps

module tfhe_pu_bd_wrapper
   (
   default_100mhz_clk_clk_n,
    default_100mhz_clk_clk_p,
    pci_express_x8_rxn,
    pci_express_x8_rxp,
    pci_express_x8_txn,
    pci_express_x8_txp,
    pcie_perstn,
    pcie_refclk_clk_n,
    pcie_refclk_clk_p,
    hbm_ref_clk_0,
    hbm_ref_clk_1,
    leds);
  input default_100mhz_clk_clk_n;
  input default_100mhz_clk_clk_p;
  input [7:0]pci_express_x8_rxn;
  input [7:0]pci_express_x8_rxp;
  output [7:0]pci_express_x8_txn;
  output [7:0]pci_express_x8_txp;
  input pcie_perstn;
  input pcie_refclk_clk_n;
  input pcie_refclk_clk_p;
  input hbm_ref_clk_0;
  input hbm_ref_clk_1;
  
  output [7:0]leds;


  wire [7:0]pci_express_x8_rxn;
  wire [7:0]pci_express_x8_rxp;
  wire [7:0]pci_express_x8_txn;
  wire [7:0]pci_express_x8_txp;
  wire pcie_perstn;
  wire pcie_refclk_clk_n;
  wire pcie_refclk_clk_p;

  tfhe_pu_bd tfhe_bd_inst
       (
       .default_100mhz_clk_clk_n(default_100mhz_clk_clk_n),
        .default_100mhz_clk_clk_p(default_100mhz_clk_clk_p),
        .pci_express_x8_rxn(pci_express_x8_rxn),
        .pci_express_x8_rxp(pci_express_x8_rxp),
        .pci_express_x8_txn(pci_express_x8_txn),
        .pci_express_x8_txp(pci_express_x8_txp),
        .pcie_perstn(pcie_perstn),
        .pcie_refclk_clk_n(pcie_refclk_clk_n),
        .pcie_refclk_clk_p(pcie_refclk_clk_p),
        .hbm_ref_clk_0(hbm_ref_clk_0),
        .hbm_ref_clk_1(hbm_ref_clk_1),
        .leds(leds)
        );
endmodule
